module alu_rol(
			input [31:0] A, B,
			output [31:0] R		//output register
);

	wire [4:0] M;			 
	assign M = B % 32;		//store modulus result in M
	//Depending on the value M rotate the 32 bit input A by B bits, bit 0 followed by bits 31 to 1 for first case
	assign R = (M == 31) ? {A[0:0], A[31:1]} :
									(M == 30) ? {A[1:0], A[31:2]} :
									(M == 29) ? {A[2:0], A[31:3]} :
												(M == 28) ? {A[3:0], A[31:4]} :
												(M == 27) ? {A[4:0], A[31:5]} :
												(M == 26) ? {A[5:0], A[31:6]} :
												(M == 25) ? {A[6:0], A[31:7]} :
												(M == 24) ? {A[7:0], A[31:8]} :
												(M == 23) ? {A[8:0], A[31:9]} :
												(M == 22) ? {A[9:0], A[31:10]} :
												(M == 21) ? {A[10:0], A[31:11]} :
												(M == 20) ? {A[11:0], A[31:12]} :
												(M == 19) ? {A[12:0], A[31:13]} :
												(M == 18) ? {A[13:0], A[31:14]} :
												(M == 17) ? {A[14:0], A[31:15]} :
												(M == 16) ? {A[15:0], A[31:16]} :
												(M == 15) ? {A[16:0], A[31:17]} :
												(M == 14) ? {A[17:0], A[31:18]} :
												(M == 13) ? {A[18:0], A[31:19]} :
												(M == 12) ? {A[19:0], A[31:20]} :
												(M == 11) ? {A[20:0], A[31:21]} :
												(M == 10) ? {A[21:0], A[31:22]} :
												(M == 9) ? {A[22:0], A[31:23]} :
												(M == 8) ? {A[23:0], A[31:24]} :
												(M == 7) ? {A[24:0], A[31:25]} :
												(M == 6) ? {A[25:0], A[31:26]} :
												(M == 5) ? {A[26:0], A[31:27]} :
												(M == 4) ? {A[27:0], A[31:28]} :
												(M == 3) ? {A[28:0], A[31:29]} :
												(M == 2) ? {A[29:0], A[31:30]} :
												(M == 1) ? {A[30:0], A[31:31]} :
												 A[31:0];
endmodule