module datapath( input R0in, R1in, R2in, R3in, R4in, R5in, R6in, R7in, R8in, R9in, R10in, R11in, R12in, R13in, R14in, R15in,
				 input R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out,
				 input wire PCin, PCout, IRin, Yin, Zin, MARin, MDRin, MDRout, HIin, HIout, LOin, LOout, IncPC, Zhighout, Zlowout, Read,
				 input AND,
				 input [31:0] MDatain,
				 input wire clk, clr
               );

                reg [15:0] enable;
                reg [15:0] Rout;

                initial begin
                    Rout = 16'b0;
                    enable = 16'b0;
                end
                
                always @* begin
                    enable[2] = R2in;
                    enable[3] = R3in;
                    enable[1] = R1in;
                    Rout[13] = R3out;
                    Rout[14] = R2out;
                end

                wire [31:0] BusMuxIn_IR, BusMuxIn_Y, C_sign_extend, BusMuxIn_InPort, BusMuxIn_MDR, BusMuxIn_PC, BusMuxIn_ZLO, BusMuxIn_ZHI, BusMuxIn_LO, BusMuxIn_HI;
                wire [31:0] BusMuxIn_R15, BusMuxIn_R14, BusMuxIn_R13, BusMuxIn_R12, BusMuxIn_R11, BusMuxIn_R10, BusMuxIn_R9, BusMuxIn_R8, BusMuxIn_R7, BusMuxIn_R6, BusMuxIn_R5, BusMuxIn_R4, BusMuxIn_R3, BusMuxIn_R2, BusMuxIn_R1, BusMuxIn_R0;
                wire [31:0] bus_signal;
                wire [31:0] C_data_out;
                wire [31:0] BusMuxOut;


                Reg32 R0(.clr(clr), .clk(clk), .Rin(enable[0]), .d(BusMuxOut), .q(busInR0));
				Reg32 R1(.clr(clr), .clk(clk), .Rin(enable[1]), .d(BusMuxOut), .q(busInR1));
				Reg32 R2(.clr(clr), .clk(clk), .Rin(enable[2]), .d(BusMuxOut), .q(busInR2));
				Reg32 R3(.clr(clr), .clk(clk), .Rin(enable[3]), .d(BusMuxOut), .q(busInR3));
				Reg32 R4(.clr(clr), .clk(clk), .Rin(enable[4]), .d(BusMuxOut), .q(busInR4));
				Reg32 R5(.clr(clr), .clk(clk), .Rin(enable[5]), .d(BusMuxOut), .q(busInR5));
				Reg32 R6(.clr(clr), .clk(clk), .Rin(enable[6]), .d(BusMuxOut), .q(busInR6));
				Reg32 R7(.clr(clr), .clk(clk), .Rin(enable[7]), .d(BusMuxOut), .q(busInR7));
				Reg32 R8(.clr(clr), .clk(clk), .Rin(enable[8]), .d(BusMuxOut), .q(busInR8));
				Reg32 R9(.clr(clr), .clk(clk), .Rin(enable[9]), .d(BusMuxOut), .q(busInR9));
				Reg32 R10(.clr(clr), .clk(clk), .Rin(enable[10]), .d(BusMuxOut), .q(busInR10));
				Reg32 R11(.clr(clr), .clk(clk), .Rin(enable[11]), .d(BusMuxOut), .q(busInR11));
				Reg32 R12(.clr(clr), .clk(clk), .Rin(enable[12]), .d(BusMuxOut), .q(busInR12));
				Reg32 R13(.clr(clr), .clk(clk), .Rin(enable[13]), .d(BusMuxOut), .q(busInR13));
				Reg32 R14(.clr(clr), .clk(clk), .Rin(enable[14]), .d(BusMuxOut), .q(busInR14));
				Reg32 R15(.clr(clr), .clk(clk), .Rin(enable[15]), .d(BusMuxOut), .q(busInR15));

                Reg32 PC(.clr(clr), .clk(clk), .Rin(PCin), .d(BusMuxOut), .q(BusMuxIn_PC));
                Reg32 Y(.clr(clr), .clk(clk), .Rin(Yin), .d(BusMuxOut), .q(BusMuxIn_Y));
                Reg32 Z_HI(.clr(clr), .clk(clk), .Rin(ZHIin), .d(C_data_out), .q(BusMuxIn_ZHI));
                Reg32 Z_LO(.clr(clr), .clk(clk), .Rin(ZLOin), .d(C_data_out), .q(BusMuxIn_ZLO));
                Reg32 HI(.clr(clr), .clk(clk), .Rin(HIin), .d(BusMuxOut), .q(BusMuxIn_HI));
                Reg32 LO(.clr(clr), .clk(clk), .Rin(LOin), .d(BusMuxOut), .q(BusMuxIn_LO));

                Reg32 IR(.clr(clr), .clk(clk), .Rin(IRin), .d(BusMuxOut), .q(BusMuxIn_IR));

                MDRreg MDR(.clr(clr), .clk(clk), .enable(MDRin), .Mdatain(Mdatain), .BusMuxOut(BusMuxOut), .Read(Read), .MDRout(BusMuxIn_MDR));

                wire[4:0] encoderOut;

                ThirtyTwoToFiveEncoder regEncoder(.Cin({{8{1'b0}},Cout,InPortout,MDRout,PCout,Zlowout,ZHighout,LOout,HIout,Rout}), .Cout(encoderOut));

                ThirtyTwoToOneEncoder busMux(
                    .BusMuxIn_R0(BusMuxIn_R0),
                    .BusMuxIn_R1(BusMuxIn_R1), 
                    .BusMuxIn_R2(BusMuxIn_R2),
                    .BusMuxIn_R3(BusMuxIn_R3),
                    .BusMuxIn_R4(BusMuxIn_R4),
                    .BusMuxIn_R5(BusMuxIn_R5),
                    .BusMuxIn_R6(BusMuxIn_R6),
                    .BusMuxIn_R7(BusMuxIn_R7),
                    .BusMuxIn_R8(BusMuxIn_R8),
                    .BusMuxIn_R9(BusMuxIn_R9),
                    .BusMuxIn_R10(BusMuxIn_R10),
                    .BusMuxIn_R11(BusMuxIn_R11),
                    .BusMuxIn_R12(BusMuxIn_R12),
                    .BusMuxIn_R13(BusMuxIn_R13),
                    .BusMuxIn_R14(BusMuxIn_R14),
                    .BusMuxIn_R15(BusMuxIn_R15),
                    .BusMuxIn_HI(BusMuxIn_HI),
                    .BusMuxIn_LO(BusMuxIn_LO),
                    .BusMuxIn_Z_high(BusMuxIn_ZHI),
                    .BusMuxIn_Z_low(BusMuxIn_ZLO),
                    .BusMuxIn_PC(BusMuxIn_PC),
                    .BusMuxIn_MDR(BusMuxIn_MDR),	
                    .BusMuxIn_InPort(BusMuxIn_InPort),
                    .C_sign_extended(C_sign_extend),
                    .BusMuxOut(BusMuxOut),
                    .select(encoderOut)
                );

                alu alu_module(
                    .Rb(BusMuxOut),
                    .Ry(BusMuxOut),
                    .AND(AND),
                    .resultLo(C_data_out)
                );


endmodule